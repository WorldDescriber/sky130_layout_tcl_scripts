magic
tech sky130A
magscale 1 2
timestamp 1771931816
<< nwell >>
rect -36 -36 234 364
rect 488 -36 758 564
<< nmos >>
rect 84 -302 114 -218
rect 608 -302 638 -134
<< pmos >>
rect 84 0 114 200
rect 608 0 638 400
<< ndiff >>
rect 524 -167 608 -134
rect 524 -201 544 -167
rect 578 -201 608 -167
rect 0 -243 84 -218
rect 0 -277 20 -243
rect 54 -277 84 -243
rect 0 -302 84 -277
rect 114 -243 198 -218
rect 114 -277 144 -243
rect 178 -277 198 -243
rect 114 -302 198 -277
rect 524 -235 608 -201
rect 524 -269 544 -235
rect 578 -269 608 -235
rect 524 -302 608 -269
rect 638 -167 722 -134
rect 638 -201 668 -167
rect 702 -201 722 -167
rect 638 -235 722 -201
rect 638 -269 668 -235
rect 702 -269 722 -235
rect 638 -302 722 -269
<< pdiff >>
rect 524 353 608 400
rect 524 319 544 353
rect 578 319 608 353
rect 524 285 608 319
rect 524 251 544 285
rect 578 251 608 285
rect 524 217 608 251
rect 0 151 84 200
rect 0 117 20 151
rect 54 117 84 151
rect 0 83 84 117
rect 0 49 20 83
rect 54 49 84 83
rect 0 0 84 49
rect 114 151 198 200
rect 114 117 144 151
rect 178 117 198 151
rect 114 83 198 117
rect 114 49 144 83
rect 178 49 198 83
rect 114 0 198 49
rect 524 183 544 217
rect 578 183 608 217
rect 524 149 608 183
rect 524 115 544 149
rect 578 115 608 149
rect 524 81 608 115
rect 524 47 544 81
rect 578 47 608 81
rect 524 0 608 47
rect 638 353 722 400
rect 638 319 668 353
rect 702 319 722 353
rect 638 285 722 319
rect 638 251 668 285
rect 702 251 722 285
rect 638 217 722 251
rect 638 183 668 217
rect 702 183 722 217
rect 638 149 722 183
rect 638 115 668 149
rect 702 115 722 149
rect 638 81 722 115
rect 638 47 668 81
rect 702 47 722 81
rect 638 0 722 47
<< ndiffc >>
rect 544 -201 578 -167
rect 20 -277 54 -243
rect 144 -277 178 -243
rect 544 -269 578 -235
rect 668 -201 702 -167
rect 668 -269 702 -235
<< pdiffc >>
rect 544 319 578 353
rect 544 251 578 285
rect 20 117 54 151
rect 20 49 54 83
rect 144 117 178 151
rect 144 49 178 83
rect 544 183 578 217
rect 544 115 578 149
rect 544 47 578 81
rect 668 319 702 353
rect 668 251 702 285
rect 668 183 702 217
rect 668 115 702 149
rect 668 47 702 81
<< psubdiff >>
rect 0 -376 198 -356
rect 0 -410 48 -376
rect 82 -410 116 -376
rect 150 -410 198 -376
rect 0 -430 198 -410
rect 524 -376 722 -356
rect 524 -410 572 -376
rect 606 -410 640 -376
rect 674 -410 722 -376
rect 524 -430 722 -410
<< nsubdiff >>
rect 524 508 722 528
rect 524 474 572 508
rect 606 474 640 508
rect 674 474 722 508
rect 524 454 722 474
rect 0 308 198 328
rect 0 274 48 308
rect 82 274 116 308
rect 150 274 198 308
rect 0 254 198 274
<< psubdiffcont >>
rect 48 -410 82 -376
rect 116 -410 150 -376
rect 572 -410 606 -376
rect 640 -410 674 -376
<< nsubdiffcont >>
rect 572 474 606 508
rect 640 474 674 508
rect 48 274 82 308
rect 116 274 150 308
<< poly >>
rect 608 400 638 430
rect 84 200 114 230
rect 84 -101 114 0
rect 356 -40 430 -20
rect 356 -74 376 -40
rect 410 -44 430 -40
rect 608 -44 638 0
rect 410 -74 638 -44
rect 356 -94 430 -74
rect 10 -121 114 -101
rect 10 -155 30 -121
rect 64 -155 114 -121
rect 608 -134 638 -74
rect 10 -175 114 -155
rect 84 -218 114 -175
rect 84 -332 114 -302
rect 608 -332 638 -302
<< polycont >>
rect 376 -74 410 -40
rect 30 -155 64 -121
<< locali >>
rect 524 508 722 524
rect 524 474 572 508
rect 606 474 640 508
rect 674 474 722 508
rect 524 458 722 474
rect 528 353 594 458
rect 528 324 544 353
rect 0 319 544 324
rect 578 319 594 353
rect 0 308 594 319
rect 0 274 48 308
rect 82 274 116 308
rect 150 285 594 308
rect 150 274 544 285
rect 0 258 544 274
rect 4 151 70 258
rect 528 251 544 258
rect 578 251 594 285
rect 528 217 594 251
rect 528 183 544 217
rect 578 183 594 217
rect 4 117 20 151
rect 54 117 70 151
rect 4 83 70 117
rect 4 49 20 83
rect 54 49 70 83
rect 4 33 70 49
rect 128 151 194 167
rect 128 117 144 151
rect 178 117 194 151
rect 128 83 194 117
rect 128 49 144 83
rect 178 49 194 83
rect 128 -27 194 49
rect 528 149 594 183
rect 528 115 544 149
rect 578 115 594 149
rect 528 81 594 115
rect 528 47 544 81
rect 578 47 594 81
rect 528 31 594 47
rect 652 353 718 369
rect 652 319 668 353
rect 702 319 718 353
rect 652 285 718 319
rect 652 251 668 285
rect 702 251 718 285
rect 652 217 718 251
rect 652 183 668 217
rect 702 183 718 217
rect 652 149 718 183
rect 652 115 668 149
rect 702 115 718 149
rect 652 81 718 115
rect 652 47 668 81
rect 702 47 718 81
rect 128 -40 426 -27
rect 128 -74 376 -40
rect 410 -74 426 -40
rect 128 -93 426 -74
rect 14 -121 80 -105
rect 14 -155 30 -121
rect 64 -155 80 -121
rect 14 -171 80 -155
rect 4 -243 70 -211
rect 4 -277 20 -243
rect 54 -277 70 -243
rect 4 -360 70 -277
rect 128 -243 194 -93
rect 128 -277 144 -243
rect 178 -277 194 -243
rect 128 -293 194 -277
rect 528 -167 594 -135
rect 528 -201 544 -167
rect 578 -201 594 -167
rect 528 -235 594 -201
rect 528 -269 544 -235
rect 578 -269 594 -235
rect 528 -360 594 -269
rect 652 -167 718 47
rect 652 -201 668 -167
rect 702 -201 718 -167
rect 652 -235 718 -201
rect 652 -269 668 -235
rect 702 -269 718 -235
rect 652 -285 718 -269
rect 0 -376 722 -360
rect 0 -410 48 -376
rect 82 -410 116 -376
rect 150 -410 572 -376
rect 606 -410 640 -376
rect 674 -410 722 -376
rect 0 -426 722 -410
<< labels >>
flabel locali 373 -77 413 -37 1 FreeSans 480 0 0 0 NET1
flabel locali 27 -158 67 -118 1 FreeSans 480 0 0 0 A
port 1 n
flabel locali 665 -272 705 -232 1 FreeSans 480 0 0 0 Y
port 2 n
flabel locali 178 271 218 311 1 FreeSans 480 0 0 0 VDD
port 3 n
flabel locali 178 -413 218 -373 1 FreeSans 480 0 0 0 VSS
port 4 n
<< end >>
