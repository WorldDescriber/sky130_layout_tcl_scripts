* NGSPICE file created from buf.ext - technology: sky130A

.subckt buf A Y VDD VSS
X0 Y.t1 NET1 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.84 pd=4.84 as=0.84 ps=4.84 w=2 l=0.15
X1 NET1 A.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.1764 pd=1.68 as=0.1764 ps=1.68 w=0.42 l=0.15
X2 Y.t0 NET1 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.3528 pd=2.52 as=0.3528 ps=2.52 w=0.84 l=0.15
X3 NET1 A.t1 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.42 pd=2.84 as=0.42 ps=2.84 w=1 l=0.15
R0 VDD.n0 VDD.t2 1243.02
R1 VDD.n1 VDD.t0 853.835
R2 VDD.n1 VDD.t1 377.945
R3 VDD.n0 VDD.t3 146.155
R4 VDD VDD.n0 70.8906
R5 VDD VDD.n1 15.1365
R6 Y.n0 Y.t1 203.329
R7 Y.n1 Y.n0 185
R8 Y.n2 Y.n1 185
R9 Y.n1 Y.t0 33.5719
R10 Y Y.n0 9.30959
R11 Y Y.n2 3.87929
R12 Y.n2 Y 3.87929
R13 A.n0 A.t1 340.089
R14 A.n0 A.t0 153.715
R15 A.n1 A.n0 152
R16 A A.n1 3.87929
R17 A.n1 A 3.87929
R18 VSS.n1 VSS.t0 737.029
R19 VSS.n1 VSS.n0 593.697
R20 VSS.n2 VSS.n1 581.737
R21 VSS.n2 VSS.t1 283.498
R22 VSS.t0 VSS.t2 232.746
R23 VSS.n0 VSS.t3 150.202
R24 VSS VSS.n0 70.4005
R25 VSS VSS.n2 15.2573
C0 A VDD 0.07328f
C1 Y VDD 0.14223f
C2 Y A 0
C3 NET1 VDD 0.20392f
C4 A NET1 0.06243f
C5 Y NET1 0.04953f
C6 Y VSS 0.21115f
C7 A VSS 0.2897f
C8 VDD VSS 1.11939f
C9 NET1 VSS 0.52746f
.ends

