** sch_path: /home/heweiwei/ask-projects/chip_project/logic_gates/not_gate/summary_working/use_sky130/inverter_2_layout_good/design_circuit/tran_inverter.sch
**.subckt tran_inverter
VIN A GND pulse(0 1.8 1n 10p 10p 5n 10n)
x1 A Y VDD GND cmos_inverter
Cload Y GND 10f m=1
VDD VDD GND 1.8
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 10p 20n
.control
run
plot V(A) V(Y)
meas tran trise TRIG V(Y) VAL=0.18 RISE=1 TARG V(Y) VAL=1.62 RISE=1
meas tran tfall TRIG V(Y) VAL=1.62 FALL=1 TARG V(Y) VAL=0.18 FALL=1
meas tran tpdr TRIG V(A) VAL=0.9 RISE=1 TARG V(Y) VAL=0.9 FALL=1
meas tran tpdf TRIG V(A) VAL=0.9 FALL=1 TARG V(Y) VAL=0.9 RISE=1
.endc


**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/heweiwei/ask-projects/chip_project/logic_gates/not_gate/summary_working/use_sky130/inverter_2_layout_good/design_circuit/inverter.sym
** sch_path: /home/heweiwei/ask-projects/chip_project/logic_gates/not_gate/summary_working/use_sky130/inverter_2_layout_good/design_circuit/inverter.sch
*.subckt inverter A Y VDD VSS
**.ipin A
**.opin Y
**.ipin VDD
**.opin VSS
*XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
*+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
*+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*.ends
.include cmos_inverter_pex.spice

.GLOBAL GND
.GLOBAL VDD
.end
