magic
tech sky130A
magscale 1 2
timestamp 1771755773
<< nwell >>
rect -36 -36 254 584
<< nmos >>
rect 94 -322 124 -122
<< pmos >>
rect 94 0 124 400
<< ndiff >>
rect 0 -171 94 -122
rect 0 -205 30 -171
rect 64 -205 94 -171
rect 0 -239 94 -205
rect 0 -273 30 -239
rect 64 -273 94 -239
rect 0 -322 94 -273
rect 124 -171 218 -122
rect 124 -205 154 -171
rect 188 -205 218 -171
rect 124 -239 218 -205
rect 124 -273 154 -239
rect 188 -273 218 -239
rect 124 -322 218 -273
<< pdiff >>
rect 0 353 94 400
rect 0 319 30 353
rect 64 319 94 353
rect 0 285 94 319
rect 0 251 30 285
rect 64 251 94 285
rect 0 217 94 251
rect 0 183 30 217
rect 64 183 94 217
rect 0 149 94 183
rect 0 115 30 149
rect 64 115 94 149
rect 0 81 94 115
rect 0 47 30 81
rect 64 47 94 81
rect 0 0 94 47
rect 124 353 218 400
rect 124 319 154 353
rect 188 319 218 353
rect 124 285 218 319
rect 124 251 154 285
rect 188 251 218 285
rect 124 217 218 251
rect 124 183 154 217
rect 188 183 218 217
rect 124 149 218 183
rect 124 115 154 149
rect 188 115 218 149
rect 124 81 218 115
rect 124 47 154 81
rect 188 47 218 81
rect 124 0 218 47
<< ndiffc >>
rect 30 -205 64 -171
rect 30 -273 64 -239
rect 154 -205 188 -171
rect 154 -273 188 -239
<< pdiffc >>
rect 30 319 64 353
rect 30 251 64 285
rect 30 183 64 217
rect 30 115 64 149
rect 30 47 64 81
rect 154 319 188 353
rect 154 251 188 285
rect 154 183 188 217
rect 154 115 188 149
rect 154 47 188 81
<< psubdiff >>
rect 0 -406 94 -376
rect 0 -440 30 -406
rect 64 -440 94 -406
rect 0 -470 94 -440
<< nsubdiff >>
rect 0 518 94 548
rect 0 484 30 518
rect 64 484 94 518
rect 0 454 94 484
<< psubdiffcont >>
rect 30 -440 64 -406
<< nsubdiffcont >>
rect 30 484 64 518
<< poly >>
rect 94 400 124 430
rect 94 -122 124 0
rect 94 -352 124 -322
<< locali >>
rect 14 518 517 534
rect 14 484 30 518
rect 64 484 517 518
rect 14 468 517 484
rect 14 353 80 468
rect 14 319 30 353
rect 64 319 80 353
rect 14 285 80 319
rect 14 251 30 285
rect 64 251 80 285
rect 14 217 80 251
rect 14 183 30 217
rect 64 183 80 217
rect 14 149 80 183
rect 14 115 30 149
rect 64 115 80 149
rect 14 81 80 115
rect 14 47 30 81
rect 64 47 80 81
rect 14 31 80 47
rect 138 353 204 369
rect 138 319 154 353
rect 188 319 204 353
rect 138 285 204 319
rect 138 251 154 285
rect 188 251 204 285
rect 138 217 204 251
rect 138 183 154 217
rect 188 183 204 217
rect 138 149 204 183
rect 138 115 154 149
rect 188 115 204 149
rect 138 81 204 115
rect 138 47 154 81
rect 188 47 204 81
rect 14 -171 80 -155
rect 14 -205 30 -171
rect 64 -205 80 -171
rect 14 -239 80 -205
rect 14 -273 30 -239
rect 64 -273 80 -239
rect 14 -390 80 -273
rect 138 -171 204 47
rect 138 -205 154 -171
rect 188 -205 204 -171
rect 138 -239 204 -205
rect 138 -273 154 -239
rect 188 -273 204 -239
rect 138 -289 204 -273
rect 14 -406 315 -390
rect 14 -440 30 -406
rect 64 -440 315 -406
rect 14 -456 315 -440
<< labels >>
flabel locali 14 468 517 534 1 FreeSans 480 0 0 0 VDD
port 3 n
flabel locali 14 -456 315 -390 1 FreeSans 480 0 0 0 VSS
port 4 n
flabel poly 94 -92 124 -30 1 FreeSans 480 0 0 0 A
port 1 n
flabel locali 138 -289 204 369 1 FreeSans 480 0 0 0 Y
port 2 n
<< end >>
