** sch_path: /home/heweiwei/ask-projects/chip_project/logic_gates/buffer_gate/use_sky130/buffer_1/design_circuit/tb_buf.sch
**.subckt tb_buf
x1 A Y VDD GND buf
Cload Y GND 10f m=1
VDD VDD GND 1.8
VA A GND pulse(0 1.8 1n 10p 10p 5n 10n)
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



* Analysis
.tran 10p 20n
.control
run
plot v(a) v(y)
* 20% to 80%
meas tran trise28 TRIG v(y) VAL=0.36 RISE=1 TARG v(y) VAL=1.44 RISE=1
* 80% to 10%
meas tran tfall82 TRIG v(y) VAL=1.44 FALL=1 TARG v(y) VAL=0.36 FALL=1
let power = v(VDD)*i(VDD)
meas tran avg_power AVG power from=1n to=20n
meas tran peak_power MAX power from=1n to=20n
meas tran trise19 TRIG V(Y) VAL=0.18 RISE=1 TARG V(Y) VAL=1.62 RISE=1
meas tran tfall91 TRIG V(Y) VAL=1.62 FALL=1 TARG V(Y) VAL=0.18 FALL=1
meas tran tpdr TRIG V(A) VAL=0.9 RISE=1 TARG V(Y) VAL=0.9 FALL=1
meas tran tpdf TRIG V(A) VAL=0.9 FALL=1 TARG V(Y) VAL=0.9 RISE=1
*(tpdr+tpdf)/2  ; Average propagation delay
meas tran energy INTEG power from=1n to=20n
*'energy/4'  ; 4 transitions in 20ns
meas tran i_peak MAX I(VDD)
meas tran i_avg AVG I(VDD) from=1n to=20n

meas tran voh MIN V(Y) from=2n to=4n   ; Output high level
meas tran vol MAX V(Y) from=7n to=9n   ; Output low level
meas tran overshoot MAX V(Y) from=1n to=3n
meas tran undershoot MIN V(Y) from=6n to=8n



.endc


***** end user architecture code
***.ends
*
** expanding   symbol:  buf.sym # of pins=4
*** sym_path: /home/heweiwei/ask-projects/chip_project/logic_gates/buffer_gate/use_sky130/buffer_1/design_circuit/buf.sym
*** sch_path: /home/heweiwei/ask-projects/chip_project/logic_gates/buffer_gate/use_sky130/buffer_1/design_circuit/buf.sch
*.subckt buf A Y VDD VSS
**.ipin A
**.opin Y
**.ipin VDD
**.ipin VSS
*x1 A net1 VDD VSS invx1
*x2 net1 Y VDD VSS invx2
*.ends
*
*
** expanding   symbol:  invx1.sym # of pins=4
*** sym_path: /home/heweiwei/ask-projects/chip_project/logic_gates/buffer_gate/use_sky130/buffer_1/design_circuit/invx1.sym
*** sch_path: /home/heweiwei/ask-projects/chip_project/logic_gates/buffer_gate/use_sky130/buffer_1/design_circuit/invx1.sch
*.subckt invx1 A Y VDD VSS
**.ipin A
**.opin Y
**.ipin VDD
**.ipin VSS
*XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
*+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
*+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*.ends
*
*
** expanding   symbol:  invx2.sym # of pins=4
*** sym_path: /home/heweiwei/ask-projects/chip_project/logic_gates/buffer_gate/use_sky130/buffer_1/design_circuit/invx2.sym
*** sch_path: /home/heweiwei/ask-projects/chip_project/logic_gates/buffer_gate/use_sky130/buffer_1/design_circuit/invx2.sch
*.subckt invx2 A Y VDD VSS
**.ipin A
**.opin Y
**.ipin VDD
**.ipin VSS
*XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
*+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
*+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
*.ends
.include buf_pex.spice

.GLOBAL GND
.GLOBAL VDD
.end
